`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//
// Create Date: 07/29/2025 08:48:20 PM
// Design Name: 
// Module Name: systolic_array_top
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module systolic_array_top #(
    parameter LEFT_MATRIX_ROW = 50,
    parameter INNER_DIMENSION = 50,
    parameter RIGHT_MATRIX_COL = 50,
    parameter DATA_WIDTH = 8 
    )(
    );
endmodule
