//////////////////////////////////////////////////////////////////////////////////
// Create Date: 01/04/2026
// Module Name: deff_vip_pkg
//////////////////////////////////////////////////////////////////////////////////

package deff_vip_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    `include "deff_vip_config.sv"
    `include "deff_vip_seq_item.sv"
    `include "deff_vip_sequencer.sv"
    `include "deff_vip_driver.sv"
    `include "deff_vip_monitor.sv"
    `include "deff_vip_agent.sv"
    `include "deff_vip_scoreboard.sv"
    `include "deff_vip_env.sv"
    `include "deff_vip_base_seq.sv"

endpackage
